module divff()
endmodule